* PEX produced on Sat Nov  9 04:40:31 AM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=2 and s=1
* NGSPICE file created from Hard_Cascode.ext - technology: sky130A

.subckt Hard_Cascode vb1 vout vinp vinn vb2 agnd avdd itail
X0 a_0_0# vb1 pfet$1_1.b agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X1 itail vinn a_1936_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X2 a_1972_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X3 vout vb2 a_1972_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=12 ps=80.6 w=40 l=0.35
X4 a_0_0# vb1 pfet$1_1.b agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4.8 ps=32.6 w=16 l=0.15
X5 a_1936_0# vb1 vout agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X6 a_1936_0# vinn itail agnd sky130_fd_pr__nfet_01v8 ad=2.4 pd=16.6 as=2 ps=8.5 w=8 l=0.15
X7 a_n436_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=6 ps=40.6 w=20 l=0.15
X8 a_n436_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X9 a_1936_0# vb1 vout agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X10 a_n436_6784# vb2 pfet$1_1.b avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X11 vout vb2 a_1972_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X12 avdd pfet$1_1.b a_1972_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X13 pfet$1_1.b vb1 a_0_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X14 avdd pfet$1_1.b a_1972_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 pfet$1_1.b vb1 a_0_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X16 vout vb1 a_1936_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X17 itail vinp a_0_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2.4 ps=16.6 w=8 l=0.15
X18 a_0_0# vinp itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X19 itail vinn a_1936_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X20 pfet$1_1.b vb2 a_n436_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X21 a_1936_0# vb1 vout agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4.8 ps=32.6 w=16 l=0.15
X22 a_1936_0# vb1 vout agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X23 itail vinp a_0_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X24 a_1936_0# vinn itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X25 pfet$1_1.b vb2 a_n436_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X26 pfet$1_1.b vb1 a_0_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4.8 pd=32.6 as=4 ps=16.5 w=16 l=0.15
X27 a_1972_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X28 vout vb2 a_1972_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X29 itail vinn a_1936_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X30 a_0_0# vinp itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X31 pfet$1_1.b vb2 a_n436_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X32 vout vb1 a_1936_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X33 a_1972_6784# vb2 vout avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X34 vout vb2 a_1972_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X35 a_0_0# vb1 pfet$1_1.b agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X36 itail vinp a_0_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X37 a_1936_0# vinn itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X38 a_n436_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X39 avdd pfet$1_1.b a_1972_6784# avdd sky130_fd_pr__pfet_01v8 ad=6 pd=40.6 as=5 ps=20.5 w=20 l=0.15
X40 a_1972_6784# vb2 vout avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X41 a_0_0# vb1 pfet$1_1.b agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X42 a_0_0# vinp itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X43 itail vinn a_1936_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X44 pfet$1_1.b vb2 a_n436_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X45 a_1936_0# vb1 vout agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X46 a_1972_6784# vb2 vout avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X47 avdd pfet$1_1.b a_n436_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X48 itail vinp a_0_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X49 a_1936_0# vinn itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X50 a_n436_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X51 itail vinp a_0_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X52 avdd pfet$1_1.b a_n436_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X53 pfet$1_1.b vb1 a_0_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X54 a_1972_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X55 a_n436_6784# vb2 pfet$1_1.b avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X56 a_0_0# vinp itail agnd sky130_fd_pr__nfet_01v8 ad=2.4 pd=16.6 as=2 ps=8.5 w=8 l=0.15
X57 a_1972_6784# vb2 vout avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X58 a_n436_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X59 a_n436_6784# vb2 pfet$1_1.b avdd sky130_fd_pr__pfet_01v8_lvt ad=12 pd=80.6 as=10 ps=40.5 w=40 l=0.35
X60 pfet$1_1.b vb2 a_n436_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=12 ps=80.6 w=40 l=0.35
X61 a_0_0# vb1 pfet$1_1.b agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X62 avdd pfet$1_1.b a_n436_6784# avdd sky130_fd_pr__pfet_01v8 ad=6 pd=40.6 as=5 ps=20.5 w=20 l=0.15
X63 avdd pfet$1_1.b a_1972_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X64 a_n436_6784# vb2 pfet$1_1.b avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X65 a_1972_6784# vb2 vout avdd sky130_fd_pr__pfet_01v8_lvt ad=12 pd=80.6 as=10 ps=40.5 w=40 l=0.35
X66 pfet$1_1.b vb1 a_0_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X67 vout vb1 a_1936_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X68 a_0_0# vinp itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
X69 avdd pfet$1_1.b a_n436_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X70 avdd pfet$1_1.b a_1972_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X71 a_n436_6784# vb2 pfet$1_1.b avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X72 itail vinn a_1936_0# agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2.4 ps=16.6 w=8 l=0.15
X73 vout vb2 a_1972_6784# avdd sky130_fd_pr__pfet_01v8_lvt ad=10 pd=40.5 as=10 ps=40.5 w=40 l=0.35
X74 vout vb1 a_1936_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4 pd=16.5 as=4 ps=16.5 w=16 l=0.15
X75 vout vb1 a_1936_0# agnd sky130_fd_pr__nfet_01v8_lvt ad=4.8 pd=32.6 as=4 ps=16.5 w=16 l=0.15
X76 avdd pfet$1_1.b a_n436_6784# avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X77 a_1972_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=6 ps=40.6 w=20 l=0.15
X78 a_1972_6784# pfet$1_1.b avdd avdd sky130_fd_pr__pfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X79 a_1936_0# vinn itail agnd sky130_fd_pr__nfet_01v8 ad=2 pd=8.5 as=2 ps=8.5 w=8 l=0.15
C0 vinn a_1936_0# 3.31006f
C1 vinp a_0_0# 3.28294f
C2 vb1 vb2 0.256342f
C3 vb2 a_1972_6784# 9.8256f
C4 avdd pfet$1_1.b 15.941099f
C5 vinp vinn 0.05232f
C6 vb1 vout 4.06787f
C7 a_n436_6784# a_1972_6784# 0.525389f
C8 vb2 a_n436_6784# 9.85438f
C9 vout a_1972_6784# 36.832897f
C10 vout vb2 9.156019f
C11 vb1 a_0_0# 3.65066f
C12 a_0_0# itail 9.55154f
C13 vb1 vinn 0.112353f
C14 vb1 a_1936_0# 3.61155f
C15 vb1 pfet$1_1.b 4.0961f
C16 vinn itail 2.92624f
C17 itail a_1936_0# 9.550059f
C18 pfet$1_1.b a_1972_6784# 3.87503f
C19 vb2 pfet$1_1.b 9.8137f
C20 vb1 avdd 0.066158f
C21 avdd a_1972_6784# 31.332802f
C22 vb1 vinp 0.112353f
C23 vb2 avdd 7.13544f
C24 a_n436_6784# pfet$1_1.b 41.466198f
C25 vout a_1936_0# 19.077599f
C26 vout pfet$1_1.b 0.257278f
C27 vinp itail 2.85599f
C28 a_n436_6784# avdd 31.3429f
C29 vout avdd 0.911318f
C30 a_0_0# a_1936_0# 0.151579f
C31 pfet$1_1.b a_0_0# 19.077599f
C32 vinn agnd 4.10322f
C33 itail agnd 4.14294f
C34 vinp agnd 4.14104f
C35 vb1 agnd 6.61838f
C36 vout agnd 7.10894f
C37 vb2 agnd 2.7681f
C38 avdd agnd 0.198677p
C39 a_1936_0# agnd 4.236701f
C40 a_0_0# agnd 4.22038f
C41 a_1972_6784# agnd 3.93674f
C42 a_n436_6784# agnd 3.91266f
C43 pfet$1_1.b agnd 12.7801f
.ends

